library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity decoder is
  port(a: in std_logic;
       b: in std_logic
)